module name();
endmodule
