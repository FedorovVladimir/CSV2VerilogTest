module NAME();
endmodule
